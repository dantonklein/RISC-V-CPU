module ram #(
    parameter int DATA_WIDTH = 32,
    parameter int ADDR_WIDTH = 32
) (

);

endmodule