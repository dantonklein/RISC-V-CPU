module branch_prediction
    
endmodule